```verilog
module TopModule(
    input logic clk,
    input logic reset,
    input logic w,
    output logic z
);

  typedef enum logic [2:0] {
    A = 3'b000,
    B = 3'b001,
    C = 3'b010,
    D = 3'b011,
    E = 3'b100,
    F = 3'b101
  } state_t;

  state_t state, next_state;

  // State transition logic
  always @(*) begin
    case (state)
      A: next_state = (w == 1'b0) ? B : A;
      B: next_state = (w == 1'b0) ? C : D;
      C: next_state = (w == 1'b0) ? E : D;
      D: next_state = (w == 1'b0) ? F : A;
      E: next_state = (w == 1'b0) ? E : D;
      F: next_state = (w == 1'b0) ? C : D;
      default: next_state = A;
    endcase
  end

  // State register
  always @(posedge clk or posedge reset) begin
    if (reset) begin
      state <= A;
    end else begin
      state <= next_state;
    end
  end

  // Output logic
  always @(*) begin
    case (state)
      E, F: z = 1'b1;
      default: z = 1'b0;
    endcase
  end

endmodule
```