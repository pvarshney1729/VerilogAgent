module TopModule (
    output logic one
);

    // Continuously drive 'one' to logic high (1)
    assign one = 1'b1;

endmodule