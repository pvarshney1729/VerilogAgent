module TopModule (
    output logic one
);

    // Always drive output one to logic high
    assign one = 1'b1;

endmodule