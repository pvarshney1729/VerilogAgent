module TopModule (
    input logic in,
    output logic out
);

    // Implementing a NOT gate
    assign out = ~in;

endmodule