module TopModule(
    output wire one
);

// Assign constant logic high to the output
assign one = 1'b1;

endmodule