```verilog
module TopModule (
  input logic in,
  output logic out
);

  // Direct combinational assignment
  assign out = in;

endmodule
```