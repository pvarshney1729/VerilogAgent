module TopModule(
    input logic in,
    output logic out
);
    // Continuous assignment for combinational logic
    assign out = in;
endmodule