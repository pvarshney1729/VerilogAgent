module TopModule (
    input  logic clk,           // Clock signal, positive edge-triggered
    input  logic areset,        // Asynchronous reset, active high
    input  logic bump_left,     // Bump from the left, active high
    input  logic bump_right,    // Bump from the right, active high
    input  logic ground,        // Ground presence, active high
    input  logic dig,           // Command to start digging, active high
    output logic walk_left,     // Lemming walking left, active high
    output logic walk_right,    // Lemming walking right, active high
    output logic aaah,          // Lemming falling, active high
    output logic digging        // Lemming digging, active high
);

    typedef enum logic [1:0] {
        STATE_WALK_LEFT = 2'b00,
        STATE_WALK_RIGHT = 2'b01,
        STATE_FALLING = 2'b10,
        STATE_DIGGING = 2'b11
    } state_t;

    state_t current_state, next_state;

    // State transition logic
    always_ff @(posedge clk or posedge areset) begin
        if (areset) begin
            current_state <= STATE_WALK_LEFT;
        end else begin
            current_state <= next_state;
        end
    end

    // Next state logic
    always_comb begin
        case (current_state)
            STATE_WALK_LEFT: begin
                if (!ground) begin
                    next_state = STATE_FALLING;
                end else if (dig) begin
                    next_state = STATE_DIGGING;
                end else if (bump_left || (bump_left && bump_right)) begin
                    next_state = STATE_WALK_RIGHT;
                end else begin
                    next_state = STATE_WALK_LEFT;
                end
            end
            STATE_WALK_RIGHT: begin
                if (!ground) begin
                    next_state = STATE_FALLING;
                end else if (dig) begin
                    next_state = STATE_DIGGING;
                end else if (bump_right) begin
                    next_state = STATE_WALK_LEFT;
                end else begin
                    next_state = STATE_WALK_RIGHT;
                end
            end
            STATE_FALLING: begin
                if (ground) begin
                    next_state = (walk_left) ? STATE_WALK_LEFT : STATE_WALK_RIGHT;
                end else begin
                    next_state = STATE_FALLING;
                end
            end
            STATE_DIGGING: begin
                if (!ground) begin
                    next_state = STATE_FALLING;
                end else begin
                    next_state = STATE_DIGGING;
                end
            end
            default: begin
                next_state = STATE_WALK_LEFT;
            end
        endcase
    end

    // Output logic
    always_comb begin
        walk_left = (current_state == STATE_WALK_LEFT);
        walk_right = (current_state == STATE_WALK_RIGHT);
        aaah = (current_state == STATE_FALLING);
        digging = (current_state == STATE_DIGGING);
    end

endmodule