module TopModule (
    input logic in,
    output logic out
);

    // Combinational logic to directly connect input to output
    assign out = in;

endmodule