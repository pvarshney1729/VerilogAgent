module TopModule(
    input  logic clk,         // Clock signal, positive edge triggered
    input  logic resetn,      // Active low synchronous reset
    input  logic x,           // Input signal from the motor
    input  logic y,           // Input signal from the motor
    output logic f,           // Output signal to control the motor
    output logic g            // Output signal to control the motor
);

    typedef enum logic [2:0] {
        STATE_A = 3'b000,
        STATE_B = 3'b001,
        STATE_C = 3'b010,
        STATE_D = 3'b011,
        STATE_E = 3'b100
    } state_t;

    state_t current_state, next_state;
    logic [1:0] x_sequence;
    logic [1:0] y_counter;

    always_ff @(posedge clk) begin
        if (!resetn) begin
            current_state <= STATE_A;
            f <= 1'b0;
            g <= 1'b0;
            x_sequence <= 2'b00;
            y_counter <= 2'b00;
        end else begin
            current_state <= next_state;
            if (current_state == STATE_B) begin
                f <= 1'b1;
            end else begin
                f <= 1'b0;
            end
            if (current_state == STATE_D) begin
                g <= 1'b1;
            end else if (current_state == STATE_E) begin
                g <= 1'b0;
            end
        end
    end

    always_comb begin
        next_state = current_state;
        case (current_state)
            STATE_A: begin
                if (resetn) begin
                    next_state = STATE_B;
                end
            end
            STATE_B: begin
                next_state = STATE_C;
            end
            STATE_C: begin
                x_sequence = {x_sequence[0], x};
                if (x_sequence == 2'b10 && x == 1'b1) begin
                    next_state = STATE_D;
                end
            end
            STATE_D: begin
                if (y == 1'b1) begin
                    next_state = STATE_D;
                end else if (y_counter == 2'b01) begin
                    next_state = STATE_E;
                end else begin
                    y_counter = y_counter + 1;
                end
            end
            STATE_E: begin
                next_state = STATE_E;
            end
            default: begin
                next_state = STATE_A;
            end
        endcase
    end

endmodule