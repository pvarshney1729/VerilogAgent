```verilog
module TopModule (
    output logic zero
);
    // Assign a constant value of 0 to the zero output
    assign zero = 1'b0;
endmodule
```