module TopModule(
    output logic output_logic_high
);

    // The combinational logic that drives the output to constant 1
    assign output_logic_high = 1'b1;

endmodule