module TopModule (
    input logic clk,           // Clock signal (1-bit, unsigned)
    input logic reset,         // Synchronous active high reset (1-bit, unsigned)
    input logic in,            // Input signal for state transitions (1-bit, unsigned)
    output logic out           // Output signal (1-bit, unsigned)
);

    // State encoding
    typedef enum logic [1:0] {
        STATE_A = 2'b00,
        STATE_B = 2'b01,
        STATE_C = 2'b10,
        STATE_D = 2'b11
    } state_t;

    state_t current_state, next_state;

    // State transition logic
    always_ff @(posedge clk) begin
        if (reset) begin
            current_state <= STATE_A;
        end else begin
            current_state <= next_state;
        end
    end

    // Next state logic
    always_comb begin
        case (current_state)
            STATE_A: begin
                if (in) 
                    next_state = STATE_B;
                else 
                    next_state = STATE_A;
            end
            STATE_B: begin
                if (in) 
                    next_state = STATE_B;
                else 
                    next_state = STATE_C;
            end
            STATE_C: begin
                if (in) 
                    next_state = STATE_D;
                else 
                    next_state = STATE_A;
            end
            STATE_D: begin
                if (in) 
                    next_state = STATE_B;
                else 
                    next_state = STATE_C;
            end
            default: next_state = STATE_A; // Default to STATE_A for safety
        endcase
    end

    // Output logic
    always_comb begin
        case (current_state)
            STATE_D: out = 1'b1;
            default: out = 1'b0;
        endcase
    end

endmodule