```verilog
module TopModule (
    output logic logic_high // Output port declaration
);

    // Constant assignment to output
    assign logic_high = 1'b1; // Drive logic high

endmodule
```