module TopModule (
    output logic out // Single-bit output, always 0
);

    // Combinational logic to drive output to 0
    assign out = 1'b0;

endmodule