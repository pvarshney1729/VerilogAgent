```verilog
module TopModule(
    output logic o_zero
);
    assign o_zero = 1'b0;
endmodule
```