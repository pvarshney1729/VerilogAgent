
// VERILOG-EVAL: response did not use [BEGIN]/[DONE] correctly