module TopModule(
    output logic zero
);
    // Assign a constant LOW (0) to the output zero
    assign zero = 1'b0;
endmodule