```verilog
[BEGIN]
module TopModule (
    input logic clk,           // Clock signal (1-bit)
    input logic reset,         // Reset signal (1-bit), active high
    input logic w,             // Input signal (1-bit)
    output logic z             // Output signal (1-bit), registered
);

// State encoding
typedef enum logic [2:0] {
    A = 3'b000,
    B = 3'b001,
    C = 3'b010,
    D = 3'b011,
    E = 3'b100,
    F = 3'b101
} state_t;

state_t current_state, next_state;

// State transition logic (combinational)
always @(*) begin
    case (current_state)
        A: next_state = (w == 1'b0) ? B : A;
        B: next_state = (w == 1'b0) ? C : D;
        C: next_state = (w == 1'b0) ? E : D;
        D: next_state = (w == 1'b0) ? F : A;
        E: next_state = (w == 1'b0) ? E : D;
        F: next_state = (w == 1'b0) ? C : D;
        default: next_state = A; // Fallback to state A
    endcase
end

// State update logic (sequential)
always @(posedge clk) begin
    if (reset) begin
        current_state <= A; // Reset to initial state A
        z <= 1'b0;          // Initialize output z
    end else begin
        current_state <= next_state; // Update state on clock edge
        z <= (current_state == E) ? 1'b1 : 1'b0; // Output logic based on state
    end
end

endmodule
[DONE]
```