module TopModule (
  input logic clk,       // Clock input, positive edge-triggered
  input logic reset,     // Reset input, synchronous active-high
  input logic w,         // 1-bit input signal
  output logic z         // 1-bit output signal
);

  typedef enum logic [2:0] {
    A = 3'b000,
    B = 3'b001,
    C = 3'b010,
    D = 3'b011,
    E = 3'b100,
    F = 3'b101
  } state_t;

  state_t current_state, next_state;

  // State transition logic
  always_ff @(posedge clk) begin
    if (reset) begin
      current_state <= A;
    end else begin
      current_state <= next_state;
    end
  end

  // Next state logic
  always_comb begin
    case (current_state)
      A: next_state = (w == 1'b0) ? B : A;
      B: next_state = (w == 1'b0) ? C : D;
      C: next_state = (w == 1'b0) ? E : D;
      D: next_state = (w == 1'b0) ? F : A;
      E: next_state = (w == 1'b0) ? E : D;
      F: next_state = (w == 1'b0) ? C : D;
      default: next_state = A; // Handle invalid states
    endcase
  end

  // Output logic
  always_comb begin
    case (current_state)
      E, F: z = 1'b1;
      default: z = 1'b0;
    endcase
  end

endmodule