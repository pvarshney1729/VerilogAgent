```verilog
module TopModule (
    input logic in,
    output logic out
);
    // Direct combinational assignment from input to output
    assign out = in;
endmodule
```