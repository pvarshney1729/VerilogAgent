module TopModule(
    input logic [7:0] a,
    input logic [7:0] b,
    input logic [7:0] c,
    input logic [7:0] d,
    output logic [7:0] min
);
    logic [7:0] min_ab, min_cd;

    assign min_ab = (a < b) ? a : b;
    assign min_cd = (c < d) ? c : d;
    assign min = (min_ab < min_cd) ? min_ab : min_cd;
endmodule