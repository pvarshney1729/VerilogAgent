module TopModule(
    input logic in,
    output logic out
);
    // Directly connect input to output
    assign out = in;
endmodule