module TopModule(
    output logic out
);

    // Drive the output 'out' to logic '0'
    assign out = 1'b0;

endmodule