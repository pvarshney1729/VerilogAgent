module TopModule(
    output logic zero
);

    // Assign zero to constant LOW
    assign zero = 1'b0;

endmodule