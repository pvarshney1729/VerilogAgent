module TopModule (
    output wire one
);
    assign one = 1'b1;
endmodule