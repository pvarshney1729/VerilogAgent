module TopModule(
    input logic in,
    output logic out
);

    // Implement NOT gate functionality
    assign out = ~in;

endmodule