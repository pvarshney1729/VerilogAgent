module TopModule (
    output logic zero // One bit output, always LOW
);

assign zero = 1'b0; // The signal 'zero' is continuously assigned to logic low (0).

endmodule