```verilog
module TopModule (
    output wire one
);
    assign one = 1'b1; // Drive the output to constant logic high
endmodule
```