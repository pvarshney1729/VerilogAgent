module TopModule (
    input logic in,
    output logic out
);
    // Direct wire connection
    assign out = in;
endmodule