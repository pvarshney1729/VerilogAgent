module TopModule (
    output logic zero
);

    // Continuous assignment to drive the output low
    assign zero = 1'b0;

endmodule