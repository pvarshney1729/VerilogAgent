module TopModule (
    input logic clk,          // Clock signal
    input logic reset,        // Active-high synchronous reset
    input logic in,           // Serial data input bit
    output logic done         // High when a valid byte is received
);

    // State encoding
    typedef enum logic [1:0] {
        IDLE = 2'b00,
        RECEIVE = 2'b01,
        VERIFY_STOP = 2'b10,
        ERROR = 2'b11
    } state_t;

    state_t current_state, next_state;
    logic [7:0] data_shift_reg;
    logic [2:0] bit_counter;

    // State transition logic
    always_ff @(posedge clk) begin
        if (reset) begin
            current_state <= IDLE;
            data_shift_reg <= 8'b0;
            bit_counter <= 3'b0;
            done <= 1'b0;
        end else begin
            current_state <= next_state;
            if (current_state == RECEIVE) begin
                data_shift_reg <= {in, data_shift_reg[7:1]};
                bit_counter <= bit_counter + 1;
            end
            if (current_state == VERIFY_STOP && in == 1'b1) begin
                done <= 1'b1;
            end else begin
                done <= 1'b0;
            end
        end
    end

    // Next state logic
    always_comb begin
        next_state = current_state;
        case (current_state)
            IDLE: begin
                if (in == 1'b0) begin
                    next_state = RECEIVE;
                end
            end
            RECEIVE: begin
                if (bit_counter == 3'b111) begin
                    next_state = VERIFY_STOP;
                end
            end
            VERIFY_STOP: begin
                if (in == 1'b1) begin
                    next_state = IDLE;
                end else begin
                    next_state = ERROR;
                end
            end
            ERROR: begin
                if (in == 1'b1) begin
                    next_state = IDLE;
                end
            end
        endcase
    end

endmodule