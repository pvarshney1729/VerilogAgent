module TopModule(
    output logic out
);
    // Assign the output to logic low (0)
    assign out = 1'b0;
endmodule