module TopModule (
    output logic out
);
    assign out = 1'b0;
endmodule