module constant_high_output(
    output logic out
);

    // Assign a constant logic high to the output
    assign out = 1'b1;

endmodule