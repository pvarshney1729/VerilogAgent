module TopModule (
    input logic in,         // 1-bit input port, unsigned
    output logic out        // 1-bit output port, unsigned
);

assign out = in;  // Direct combinational assignment

endmodule