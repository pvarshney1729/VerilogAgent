module TopModule(
    input [254:0] in_vector,
    output [7:0] out_count
);

    assign out_count = in_vector[0] + in_vector[1] + in_vector[2] + in_vector[3] +
                       in_vector[4] + in_vector[5] + in_vector[6] + in_vector[7] +
                       in_vector[8] + in_vector[9] + in_vector[10] + in_vector[11] +
                       in_vector[12] + in_vector[13] + in_vector[14] + in_vector[15] +
                       in_vector[16] + in_vector[17] + in_vector[18] + in_vector[19] +
                       in_vector[20] + in_vector[21] + in_vector[22] + in_vector[23] +
                       in_vector[24] + in_vector[25] + in_vector[26] + in_vector[27] +
                       in_vector[28] + in_vector[29] + in_vector[30] + in_vector[31] +
                       in_vector[32] + in_vector[33] + in_vector[34] + in_vector[35] +
                       in_vector[36] + in_vector[37] + in_vector[38] + in_vector[39] +
                       in_vector[40] + in_vector[41] + in_vector[42] + in_vector[43] +
                       in_vector[44] + in_vector[45] + in_vector[46] + in_vector[47] +
                       in_vector[48] + in_vector[49] + in_vector[50] + in_vector[51] +
                       in_vector[52] + in_vector[53] + in_vector[54] + in_vector[55] +
                       in_vector[56] + in_vector[57] + in_vector[58] + in_vector[59] +
                       in_vector[60] + in_vector[61] + in_vector[62] + in_vector[63] +
                       in_vector[64] + in_vector[65] + in_vector[66] + in_vector[67] +
                       in_vector[68] + in_vector[69] + in_vector[70] + in_vector[71] +
                       in_vector[72] + in_vector[73] + in_vector[74] + in_vector[75] +
                       in_vector[76] + in_vector[77] + in_vector[78] + in_vector[79] +
                       in_vector[80] + in_vector[81] + in_vector[82] + in_vector[83] +
                       in_vector[84] + in_vector[85] + in_vector[86] + in_vector[87] +
                       in_vector[88] + in_vector[89] + in_vector[90] + in_vector[91] +
                       in_vector[92] + in_vector[93] + in_vector[94] + in_vector[95] +
                       in_vector[96] + in_vector[97] + in_vector[98] + in_vector[99] +
                       in_vector[100] + in_vector[101] + in_vector[102] + in_vector[103] +
                       in_vector[104] + in_vector[105] + in_vector[106] + in_vector[107] +
                       in_vector[108] + in_vector[109] + in_vector[110] + in_vector[111] +
                       in_vector[112] + in_vector[113] + in_vector[114] + in_vector[115] +
                       in_vector[116] + in_vector[117] + in_vector[118] + in_vector[119] +
                       in_vector[120] + in_vector[121] + in_vector[122] + in_vector[123] +
                       in_vector[124] + in_vector[125] + in_vector[126] + in_vector[127] +
                       in_vector[128] + in_vector[129] + in_vector[130] + in_vector[131] +
                       in_vector[132] + in_vector[133] + in_vector[134] + in_vector[135] +
                       in_vector[136] + in_vector[137] + in_vector[138] + in_vector[139] +
                       in_vector[140] + in_vector[141] + in_vector[142] + in_vector[143] +
                       in_vector[144] + in_vector[145] + in_vector[146] + in_vector[147] +
                       in_vector[148] + in_vector[149] + in_vector[150] + in_vector[151] +
                       in_vector[152] + in_vector[153] + in_vector[154] + in_vector[155] +
                       in_vector[156] + in_vector[157] + in_vector[158] + in_vector[159] +
                       in_vector[160] + in_vector[161] + in_vector[162] + in_vector[163] +
                       in_vector[164] + in_vector[165] + in_vector[166] + in_vector[167] +
                       in_vector[168] + in_vector[169] + in_vector[170] + in_vector[171] +
                       in_vector[172] + in_vector[173] + in_vector[174] + in_vector[175] +
                       in_vector[176] + in_vector[177] + in_vector[178] + in_vector[179] +
                       in_vector[180] + in_vector[181] + in_vector[182] + in_vector[183] +
                       in_vector[184] + in_vector[185] + in_vector[186] + in_vector[187] +
                       in_vector[188] + in_vector[189] + in_vector[190] + in_vector[191] +
                       in_vector[192] + in_vector[193] + in_vector[194] + in_vector[195] +
                       in_vector[196] + in_vector[197] + in_vector[198] + in_vector[199] +
                       in_vector[200] + in_vector[201] + in_vector[202] + in_vector[203] +
                       in_vector[204] + in_vector[205] + in_vector[206] + in_vector[207] +
                       in_vector[208] + in_vector[209] + in_vector[210] + in_vector[211] +
                       in_vector[212] + in_vector[213] + in_vector[214] + in_vector[215] +
                       in_vector[216] + in_vector[217] + in_vector[218] + in_vector[219] +
                       in_vector[220] + in_vector[221] + in_vector[222] + in_vector[223] +
                       in_vector[224] + in_vector[225] + in_vector[226] + in_vector[227] +
                       in_vector[228] + in_vector[229] + in_vector[230] + in_vector[231] +
                       in_vector[232] + in_vector[233] + in_vector[234] + in_vector[235] +
                       in_vector[236] + in_vector[237] + in_vector[238] + in_vector[239] +
                       in_vector[240] + in_vector[241] + in_vector[242] + in_vector[243] +
                       in_vector[244] + in_vector[245] + in_vector[246] + in_vector[247] +
                       in_vector[248] + in_vector[249] + in_vector[250] + in_vector[251] +
                       in_vector[252] + in_vector[253] + in_vector[254];

endmodule