module TopModule(
    output logic one
);

    // Assign the constant value 1 to the output 'one'
    assign one = 1'b1;

endmodule