module TopModule
(
  output logic one
);

  // Combinational logic

  assign one = 1'b1;

endmodule