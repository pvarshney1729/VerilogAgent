module TopModule (
    input logic in_signal,
    output logic out_signal
);

    assign out_signal = in_signal;

endmodule