module TopModule(
    input logic in,
    output logic out
);
    // Implementing NOT gate
    assign out = ~in;
endmodule