```verilog
[BEGIN]
module TopModule (
    input logic clk,           // Clock signal (rising edge triggered)
    input logic load,         // Load signal (active high)
    input logic ena,          // Enable signal for shifting (active high)
    input logic [1:0] amount, // Shift amount control
    input logic [63:0] data,  // Data to load into the shift register (unsigned 64-bit)
    output logic [63:0] q     // Shift register output (unsigned 64-bit)
);

always @(posedge clk) begin
    if (load) begin
        q <= data; // Load data into shift register
    end else if (ena) begin
        case (amount)
            2'b00: q <= {q[62:0], 1'b0}; // Shift left by 1 bit
            2'b01: q <= {q[55:0], 8'b0}; // Shift left by 8 bits
            2'b10: q <= {q[63], q[62:1]}; // Arithmetic shift right by 1 bit
            2'b11: q <= {q[63], q[63:8]}; // Arithmetic shift right by 8 bits
        endcase
    end
end

endmodule
[DONE]
```