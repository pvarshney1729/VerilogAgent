module TopModule (
    input logic in,
    output logic out
);

    // Assign the output to the same value as the input
    assign out = in;

endmodule