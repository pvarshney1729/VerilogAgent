module TopModule(
    output logic zero
);

    // Assign zero to always output LOW
    assign zero = 1'b0;

endmodule