```verilog
module TopModule(
    output logic one
);

// Assign constant logic high to the output
assign one = 1'b1;

endmodule
```