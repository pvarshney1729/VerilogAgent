module TopModule
(
  output logic zero
);

  // Combinational logic

  assign zero = 0;

endmodule