module TopModule (
    output logic out
);
    // Combinational assignment
    assign out = 1'b0;
endmodule