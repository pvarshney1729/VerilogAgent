module TopModule(
    output logic out
);

    // Drive the output 'out' to logic low (0)
    assign out = 1'b0;

endmodule