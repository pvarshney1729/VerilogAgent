```
[BEGIN]
module TopModule (
    input logic clk,
    input logic reset,
    output logic [2:0] ena,
    output logic [15:0] q
);
    always @(posedge clk) begin
        if (reset) begin
            q <= 16'b0000_0000_0000_0000;
            ena <= 3'b000;
        end else begin
            ena <= 3'b000; // Clear enable signals
            
            // Increment Ones Digit
            if (q[3:0] == 4'd9) begin
                q[3:0] <= 4'b0000;
                ena[0] <= 1'b1; // Enable for ones digit
                // Increment Tens Digit
                if (q[7:4] == 4'd9) begin
                    q[7:4] <= 4'b0000;
                    ena[1] <= 1'b1; // Enable for tens digit
                    // Increment Hundreds Digit
                    if (q[11:8] == 4'd9) begin
                        q[11:8] <= 4'b0000;
                        ena[2] <= 1'b1; // Enable for hundreds digit
                        // Increment Thousands Digit
                        if (q[15:12] == 4'd9) begin
                            q <= 16'b0000_0000_0000_0000; // Reset to 0
                        end else begin
                            q[15:12] <= q[15:12] + 1'b1;
                        end
                    end else begin
                        q[11:8] <= q[11:8] + 1'b1;
                    end
                end else begin
                    q[7:4] <= q[7:4] + 1'b1;
                end
            end else begin
                q[3:0] <= q[3:0] + 1'b1;
            end
        end
    end
endmodule
[DONE]
```