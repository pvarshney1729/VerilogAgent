```verilog
[BEGIN]
module TopModule (
    input logic clk,
    input logic reset,
    input logic j,
    input logic k,
    output logic out
);

    // State encoding
    localparam logic OFF = 1'b0;
    localparam logic ON  = 1'b1;
    
    // State registers
    logic state, next_state;

    // State transition logic
    always @(posedge clk) begin
        if (reset) begin
            state <= OFF;
        end else begin
            state <= next_state;
        end
    end

    // Next state logic
    always @(*) begin
        case (state)
            OFF: begin
                if (j)
                    next_state = ON;
                else
                    next_state = OFF;
            end
            ON: begin
                if (k)
                    next_state = OFF;
                else
                    next_state = ON;
            end
            default: next_state = OFF;
        endcase
    end

    // Output logic
    always @(*) begin
        out = (state == ON) ? 1'b1 : 1'b0;
    end

endmodule
[DONE]
```