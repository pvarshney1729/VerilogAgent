module TopModule (
    input logic [2:0] y,
    input logic w,
    input logic clk,
    input logic reset,
    output logic Y1
);

    logic [2:0] state, next_state;

    // State transition logic
    always @(*) begin
        case (state)
            3'b000: next_state = (w == 0) ? 3'b001 : 3'b000; // State A
            3'b001: next_state = (w == 0) ? 3'b010 : 3'b011; // State B
            3'b010: next_state = (w == 0) ? 3'b100 : 3'b011; // State C
            3'b011: next_state = (w == 0) ? 3'b101 : 3'b000; // State D
            3'b100: next_state = (w == 0) ? 3'b100 : 3'b011; // State E
            3'b101: next_state = (w == 0) ? 3'b010 : 3'b011; // State F
            default: next_state = 3'b000; // Undefined states transition to State A
        endcase
    end

    // State register with asynchronous reset
    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            state <= 3'b000; // Initialize to State A
        end else begin
            state <= next_state;
        end
    end

    // Output logic
    assign Y1 = state[1];

endmodule