module TopModule
(
  input  logic in,
  output logic out
);

  // Combinational logic

  assign out = ~in;

endmodule