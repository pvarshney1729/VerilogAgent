```verilog
module TopModule(
    output logic logic_high
);
    // Drive logic high (1) on the output
    assign logic_high = 1'b1;
endmodule
```