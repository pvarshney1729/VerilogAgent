module TopModule (
    input  logic [3:0] x,
    output logic f
);
    assign f = (x[3:2] == 2'b11 && x[1:0] == 2'b00) || // 1 (11, 00)
               (x[3:2] == 2'b11 && x[1:0] == 2'b01) || // 1 (11, 01)
               (x[3:2] == 2'b01 && x[1:0] == 2'b10) || // 1 (01, 10)
               (x[3:2] == 2'b10 && x[1:0] == 2'b00) || // 1 (10, 00)
               (x[3:2] == 2'b10 && x[1:0] == 2'b01);   // 1 (10, 01)
endmodule