module TopModule (
    output logic high_signal
);

    // Continuous assignment to drive the output high
    assign high_signal = 1'b1;

endmodule