module top_module (
    output logic zero  // 1-bit combinational output, always LOW
);

// Assign a constant logic LOW to the output
assign zero = 1'b0;

endmodule