module TopModule (
    output logic out_zero // Clarified output name and type
);

    // Combinational assignment
    assign out_zero = 1'b0; // Explicitly specify the bit width and value

endmodule