```verilog
module TopModule(
  output logic out  // Define the output as a single-bit logic type 
);
  // Assign a constant value of 0 to the output
  assign out = 1'b0;  // Explicitly indicate a 1-bit binary constant

endmodule
```