```verilog
module TopModule (
    output logic out // Define the output as logic
);

    // Assign the output to logic low
    assign out = 1'b0;

endmodule
```