module TopModule (
    output wire out
);
    // Continuous assignment to drive 'out' to logic low
    assign out = 1'b0;
endmodule