module TopModule (
    output logic out
);
    assign out = 1'b0; // Drive out to logic low (0) continuously
endmodule