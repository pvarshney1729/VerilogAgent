module TopModule (
    input  logic a,
    input  logic b,
    input  logic cin,
    output logic cout,
    output logic sum
);

    always @(*) begin
        // Full adder logic
        sum  = a ^ b ^ cin;
        cout = (a & b) | (b & cin) | (cin & a);
    end

endmodule