module TopModule (
    output wire zero  // Single-bit output port named 'zero'
);

    // Assign constant logic LOW to the output 'zero'
    assign zero = 1'b0;

endmodule