module TopModule (
    input wire a,
    input wire b,
    input wire c,
    input wire d,
    output wire out,
    output wire out_n
);

    // Internal wire declarations
    wire and1_out;
    wire and2_out;

    // AND gate logic
    assign and1_out = a & b;
    assign and2_out = c & d;

    // OR gate logic
    assign out = and1_out | and2_out;

    // NOT gate logic
    assign out_n = ~out;

endmodule