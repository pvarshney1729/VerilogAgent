module TopModule (
    output logic out
);

    // Continuous assignment to drive output to 0
    assign out = 1'b0;

endmodule