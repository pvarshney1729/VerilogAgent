module TopModule (
    output logic out // Output port named 'out' of type logic; 1-bit width
);

assign out = 1'b1; // Assign logic high to the output

endmodule