module TopModule (
    input  logic clk,
    input  logic areset,
    input  logic [7:0] d,
    output logic [7:0] q
);

    always @(posedge clk or posedge areset) begin
        if (areset) begin
            q <= 8'b00000000; // Reset all outputs to 0
        end else begin
            q <= d; // Capture input d on the positive edge of clk
        end
    end

endmodule