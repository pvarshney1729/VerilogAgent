module TopModule (
    logic a,
    logic b,
    logic out
);
    // AND gate implementation
    assign out = a & b;
endmodule