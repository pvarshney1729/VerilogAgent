module TopModule(
    output logic one
);

    // Assign a constant logic high to the output
    assign one = 1'b1;

endmodule