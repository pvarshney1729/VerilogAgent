module TopModule
(
  output logic out
);

  // Combinational logic

  assign out = 0;

endmodule