[BEGIN]
module TopModule (
    output logic out  // Use 'logic' type for output
);

// Assign a constant logic low (0) directly to the output 'out'
assign out = 1'b0;

endmodule
[DONE]