module TopModule(
    input wire in,
    output wire out
);
    // Directly connect the input to the output
    assign out = in;
endmodule