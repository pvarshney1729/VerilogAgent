module TopModule(
    input logic a,
    input logic b,
    output logic q
);
    // Implementing the AND operation
    assign q = a & b;
endmodule