```verilog
module TopModule (
    input logic in,
    output logic out
);
    // Direct assignment to mimic wire behavior
    assign out = in;
endmodule
```