module TopModule(
    input logic clk,
    input logic reset,
    output logic [3:0] q
);

    // Initial state for simulation
    initial begin
        q = 4'b0000;
    end

    // Sequential logic for counter with synchronous reset
    always_ff @(posedge clk) begin
        if (reset) begin
            q <= 4'b0000;
        end else begin
            q <= q + 1'b1;
        end
    end

endmodule