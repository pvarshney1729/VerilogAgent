module TopModule (
    input logic [3:0] x,  // x[3] (MSB), x[2], x[1], x[0] (LSB)
    output logic f        // 1-bit output
);

    assign f = (x[3] & ~x[2] & ~x[1] & x[0]) | 
               (~x[3] & x[2] & x[1]) | 
               (x[3] & x[2] & ~x[1] & x[0]) | 
               (x[2] & ~x[3] & x[1] & x[0]);

endmodule