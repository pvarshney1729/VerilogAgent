module TopModule(
  output logic one
);
  assign one = 1'b1; // Drive the output to logic high
endmodule