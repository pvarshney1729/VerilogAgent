module TopModule
(
  input  logic [3:0] a,
  input  logic [3:0] b,
  input  logic [3:0] c,
  input  logic [3:0] d,
  input  logic [3:0] e,
  output logic [3:0] q
);

  // Combinational logic

  always @(*) begin
    case (c)
      4'b0000: q = b;
      4'b0001: q = e;
      4'b0010: q = a;
      4'b0011: q = d;
      default:  q = 4'b1111;
    endcase
  end

endmodule