```verilog
module pattern_detector (
    input logic clk,
    input logic reset,
    input logic data_in,
    output logic pattern_detected
);

    typedef enum logic [2:0] {
        IDLE = 3'b000,
        S1   = 3'b001,
        S11  = 3'b010,
        S110 = 3'b011,
        S1101= 3'b100
    } state_t;

    state_t current_state, next_state;

    // State transition logic
    always_ff @(posedge clk) begin
        if (reset) begin
            current_state <= IDLE;
        end else begin
            current_state <= next_state;
        end
    end

    // Next state logic
    always @(*) begin
        case (current_state)
            IDLE:  next_state = (data_in) ? S1 : IDLE;
            S1:    next_state = (data_in) ? S11 : IDLE;
            S11:   next_state = (data_in) ? S11 : S110;
            S110:  next_state = (data_in) ? S1101 : IDLE;
            S1101: next_state = (data_in) ? S11 : IDLE;
            default: next_state = IDLE;
        endcase
    end

    // Output logic
    always @(*) begin
        pattern_detected = (current_state == S1101);
    end

endmodule
```