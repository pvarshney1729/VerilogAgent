module TopModule(
    input  logic in,
    output logic out
);

    // Combinational assignment
    assign out = in;

endmodule