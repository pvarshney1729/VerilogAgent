module TopModule (
    input logic x,
    input logic y,
    output logic z
);

    // Implement the boolean function z = (x^y) & x
    always @(*) begin
        z = (x ^ y) & x;
    end

endmodule