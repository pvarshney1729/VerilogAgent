module TopModule (
    output logic out
);
    // Constantly drive output to logic low
    assign out = 1'b0;
endmodule