module TopModule (
    output logic zero
);

    assign zero = 1'b0; // Continuously drive output 'zero' to LOW

endmodule