```verilog
module TopModule (
    output logic zero
);

// Assign the output to a constant LOW
assign zero = 1'b0;

endmodule
```