module TopModule (
    input logic in,
    output logic out
);

    // Directly propagate the input to the output
    assign out = in;

endmodule