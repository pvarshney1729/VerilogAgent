module TopModule(
    input [3:0] x,
    output logic f
);

always @(*) begin
    case (x)
        4'b0101, 4'b0110, 4'b1000, 4'b1001, 4'b1100, 4'b1101, 4'b1110: f = 1'b1;
        4'b0001, 4'b0010, 4'b0100: f = 1'b0;
        default: f = 1'bx; // Don't-care conditions
    endcase
end

endmodule