module TopModule (
    input  logic in,
    output logic out
);

    // Implement NOT gate using assign statement
    assign out = ~in;

endmodule