```
[BEGIN]
module TopModule (
    output logic zero
);
    // Constantly assign zero to the output
    assign zero = 1'b0;
endmodule
[DONE]
```