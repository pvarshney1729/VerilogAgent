```verilog
module TopModule (
    output logic one
);

// Continuous assignment to drive the output high
assign one = 1'b1;

endmodule
```