module TopModule (
    output logic zero
);

// Constantly drive `zero` to 0
assign zero = 1'b0;

endmodule