module TopModule (
    output logic out
);

    // Always drive out to logic low
    assign out = 1'b0;

endmodule