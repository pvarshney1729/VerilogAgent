module TopModule (
    input logic in_bit,   // Single-bit input signal
    output logic out_bit  // Single-bit output signal
);

    assign out_bit = in_bit; // Combinational assignment

endmodule