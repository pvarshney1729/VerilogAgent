```verilog
module TopModule (
    output logic out
);
    // Assign the output to logic low
    assign out = 1'b0;
endmodule
```