module TopModule(
    input logic in,
    output logic out
);
    // Implementing NOT gate logic
    assign out = ~in;
endmodule