module TopModule(
    output logic one
);
    // Constantly drive the output high
    assign one = 1'b1;
endmodule