module TopModule (
    logic in,
    logic out
);
    assign out = ~in;
endmodule