module TopModule(
    output logic logic_high
);

    // Constantly drive the output to logic high
    assign logic_high = 1'b1;

endmodule