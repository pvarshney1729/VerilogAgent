module TopModule(
    output logic zero
);
    // Continuous assignment to set the output 'zero' to logical LOW
    assign zero = 1'b0;
endmodule