module WireModule(
    input logic in,      // One-bit input signal
    output logic out     // One-bit output signal
);

assign out = in; // Direct connection

endmodule