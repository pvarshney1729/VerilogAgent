module TopModule (
    output logic zero
);
    // Continuous assignment to drive output zero to logic LOW
    assign zero = 1'b0;

endmodule