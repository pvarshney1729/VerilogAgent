module TopModule(
    output logic out
);
    // Constant drive of logic low
    assign out = 1'b0;
endmodule