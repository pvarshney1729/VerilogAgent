module TopModule (
    logic a,
    logic b,
    logic c,
    logic out
);
    // Implementing the simplified logic derived from the Karnaugh map
    assign out = b;
endmodule