module TopModule (
    input logic clk,
    input logic reset,
    input logic data,
    output logic start_shifting
);
    typedef enum logic [2:0] {
        S0, // Initial state
        S1, // Received 1
        S2, // Received 11
        S3  // Received 110
    } state_t;

    state_t current_state, next_state;

    always_ff @(posedge clk) begin
        if (reset) begin
            current_state <= S0;
            start_shifting <= 1'b0;
        end else begin
            current_state <= next_state;
        end
    end

    always_ff @(posedge clk) begin
        if (reset) begin
            start_shifting <= 1'b0;
        end else if (current_state == S3 && data == 1'b1) begin
            start_shifting <= 1'b1;
        end
    end

    always_comb begin
        case (current_state)
            S0: begin
                if (data == 1'b1) 
                    next_state = S1;
                else 
                    next_state = S0;
            end
            S1: begin
                if (data == 1'b1) 
                    next_state = S2;
                else 
                    next_state = S0;
            end
            S2: begin
                if (data == 1'b0) 
                    next_state = S3;
                else 
                    next_state = S2;
            end
            S3: begin
                if (data == 1'b1) 
                    next_state = S1;
                else 
                    next_state = S0;
            end
            default: next_state = S0;
        endcase
    end
endmodule