module TopModule(
    output logic one
);
    assign one = 1'b1; // Always drive the output to logic high
endmodule