module TopModule(
    output logic one
);

    // Drive the output 'one' to logic high
    assign one = 1'b1;

endmodule