module TopModule (
    output logic out
);

    assign out = 1'b0; // Always drive output to logic low

endmodule