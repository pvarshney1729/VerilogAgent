module TopModule(
    output logic out
);
    // Assign a constant logic low to the output
    assign out = 1'b0;
endmodule