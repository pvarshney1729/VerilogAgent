```verilog
module TopModule (
    input logic in,  // Single-bit input signal
    output logic out // Single-bit output signal
);

// Combinational assignment
assign out = in;

endmodule
```