module TopModule (
    input logic clk,
    input logic rst,
    input logic shift_ena,
    input logic count_ena,
    input logic data,
    output logic [3:0] q
);

    always_ff @(posedge clk) begin
        if (rst) begin
            q <= 4'b0000;
        end else if (shift_ena && !count_ena) begin
            q <= {q[2:0], data};
        end else if (count_ena && !shift_ena) begin
            q <= q - 1'b1;
        end
        // Undefined behavior if both shift_ena and count_ena are high
    end

endmodule