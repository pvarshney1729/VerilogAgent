module TopModule (
    input  logic clk,
    input  logic reset,
    input  logic in,
    output logic disc,
    output logic flag,
    output logic err
);

    typedef enum logic [2:0] {
        S0, // Initial state
        S1, // Received 1
        S2, // Received 11
        S3, // Received 111
        S4, // Received 1111
        S5, // Received 11111
        S6, // Received 111111
        S7  // Received 1111111 (error state)
    } state_t;

    state_t state, next_state;

    // Sequential logic for state transition
    always @(posedge clk) begin
        if (reset) begin
            state <= S0;
        end else begin
            state <= next_state;
        end
    end

    // Combinational logic for next state and outputs
    always @(*) begin
        next_state = state;
        disc = 1'b0;
        flag = 1'b0;
        err = 1'b0;

        case (state)
            S0: begin
                if (in) next_state = S1;
            end
            S1: begin
                if (in) next_state = S2;
                else next_state = S0;
            end
            S2: begin
                if (in) next_state = S3;
                else next_state = S0;
            end
            S3: begin
                if (in) next_state = S4;
                else next_state = S0;
            end
            S4: begin
                if (in) next_state = S5;
                else next_state = S0;
            end
            S5: begin
                if (in) next_state = S6;
                else next_state = S0;
            end
            S6: begin
                if (in) begin
                    next_state = S7; // Error state
                    err = 1'b1; // Signal error
                end else begin
                    next_state = S0; // Reset to initial state
                    disc = 1'b1; // Signal discard
                end
            end
            S7: begin
                // Stay in error state
                err = 1'b1; // Signal error
                if (!in) next_state = S0; // Reset to initial state on 0
            end
        endcase

        // Flag output for frame boundaries
        if (state == S6 && in) begin
            flag = 1'b1; // Signal flag
        end
    end

endmodule