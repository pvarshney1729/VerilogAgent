module TopModule(
    input  logic in,
    output logic out
);

    // Combinational logic to assign the output to the input
    assign out = in;

endmodule