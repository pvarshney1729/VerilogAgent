module TopModule(
    output logic out
);

    // Assign a constant value of 0 to the output
    assign out = 1'b0;

endmodule