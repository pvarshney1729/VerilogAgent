module TopModule (
    input logic clk,
    input logic reset,
    input logic s,
    input logic w,
    output logic z
);

    typedef enum logic [1:0] {
        STATE_A = 2'b00,
        STATE_B = 2'b01
    } state_t;

    state_t current_state, next_state;
    logic [1:0] w_counter;
    logic [1:0] cycle_counter;

    always_ff @(posedge clk) begin
        if (reset) begin
            current_state <= STATE_A;
            w_counter <= 2'b00;
            cycle_counter <= 2'b00;
            z <= 1'b0;
        end else begin
            current_state <= next_state;
            if (current_state == STATE_B) begin
                cycle_counter <= cycle_counter + 1;
                if (w) begin
                    w_counter <= w_counter + 1;
                end
                if (cycle_counter == 2'b10) begin
                    z <= (w_counter == 2'b10) ? 1'b1 : 1'b0;
                    w_counter <= 2'b00;
                    cycle_counter <= 2'b00;
                end
            end
        end
    end

    always_comb begin
        case (current_state)
            STATE_A: begin
                if (s) begin
                    next_state = STATE_B;
                end else begin
                    next_state = STATE_A;
                end
            end
            STATE_B: begin
                next_state = STATE_B;
            end
            default: begin
                next_state = STATE_A;
            end
        endcase
    end

endmodule