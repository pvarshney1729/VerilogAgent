module TopModule(
    input logic in,
    output logic out
);

    // Combinational logic to assign output to input
    assign out = in;

endmodule