```verilog
module TopModule (
    input logic in,
    output logic out
);
    // Combinational assignment of output to input
    assign out = in;
endmodule
```