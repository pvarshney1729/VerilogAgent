module TopModule(
    output logic zero
);

    // Assign the output 'zero' to a constant LOW
    assign zero = 1'b0;

endmodule