module TopModule (
    input logic i_in,
    output logic o_out
);

    // Combinational logic: direct assignment
    assign o_out = i_in;

endmodule