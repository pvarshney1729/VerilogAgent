module TopModule (
    input  logic p1a,  // 1-bit input
    input  logic p1b,  // 1-bit input
    input  logic p1c,  // 1-bit input
    input  logic p1d,  // 1-bit input
    input  logic p1e,  // 1-bit input
    input  logic p1f,  // 1-bit input
    input  logic p2a,  // 1-bit input
    input  logic p2b,  // 1-bit input
    input  logic p2c,  // 1-bit input
    input  logic p2d,  // 1-bit input
    output logic p1y,  // 1-bit output
    output logic p2y   // 1-bit output
);

    logic and1_out, and2_out, and3_out, and4_out;

    assign and1_out = p1a & p1b & p1c;
    assign and2_out = p1d & p1e & p1f;
    assign and3_out = p2a & p2b;
    assign and4_out = p2c & p2d;

    assign p1y = and1_out | and2_out;
    assign p2y = and3_out | and4_out;

endmodule