module TopModule (
    input wire in,    // 1-bit unsigned input
    output wire out   // 1-bit unsigned output
);
    // Combinational logic: direct assignment
    assign out = in;

endmodule