module AndGate (
    input wire a,
    input wire b,
    output wire q
);

assign q = a & b;

endmodule