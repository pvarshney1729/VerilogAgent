module TopModule (
    input logic clk,               // Clock signal, active on positive edge
    input logic reset,             // Active-high synchronous reset
    input logic data,              // Data input stream, 1-bit wide
    output logic start_shifting     // Output signal, set to 1 when sequence is found
);

    typedef enum logic [2:0] {
        IDLE = 3'b000,
        S1   = 3'b001,
        S11  = 3'b010,
        S110 = 3'b011,
        MATCHED = 3'b100
    } state_t;

    state_t current_state, next_state;

    always_ff @(posedge clk) begin
        if (reset) begin
            current_state <= IDLE;
            start_shifting <= 1'b0;
        end else begin
            current_state <= next_state;
        end
    end

    always_comb begin
        case (current_state)
            IDLE: begin
                if (data) begin
                    next_state = S1;
                end else begin
                    next_state = IDLE;
                end
                start_shifting = 1'b0;
            end
            S1: begin
                if (data) begin
                    next_state = S11;
                end else begin
                    next_state = IDLE;
                end
                start_shifting = 1'b0;
            end
            S11: begin
                if (data) begin
                    next_state = S110;
                end else begin
                    next_state = IDLE;
                end
                start_shifting = 1'b0;
            end
            S110: begin
                if (!data) begin
                    next_state = MATCHED;
                end else begin
                    next_state = S11;
                end
                start_shifting = 1'b0;
            end
            MATCHED: begin
                start_shifting = 1'b1;
                next_state = IDLE; // or remain in MATCHED based on further requirements
            end
            default: begin
                next_state = IDLE;
                start_shifting = 1'b0;
            end
        endcase
    end

endmodule