```verilog
[BEGIN]
module TopModule (
    output logic zero
);
    always @(*) begin
        zero = 1'b0;
    end
endmodule
[DONE]
```