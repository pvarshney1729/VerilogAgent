module TopModule (
    output logic output_one
);

    // Continuously drive the output to logic high
    assign output_one = 1'b1;

endmodule