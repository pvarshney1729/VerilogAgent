module TopModule(output logic zero);
  assign zero = 1'b0;
endmodule