module TopModule(
    output logic out
);

    // Always drive the output to 0
    assign out = 1'b0;

endmodule