module TopModule (
    input logic clk,  // Clock signal, positive edge-triggered
    input logic x,    // Single-bit input
    output logic z    // Single-bit output
);

    logic dff1, dff2, dff3;
    logic xor_out, and_out, or_out;

    // Combinational logic for gates
    always @(*) begin
        xor_out = x ^ dff1;
        and_out = x & ~dff2;
        or_out  = x | ~dff3;
    end

    // Sequential logic for D flip-flops with asynchronous reset
    always_ff @(posedge clk) begin
        dff1 <= xor_out;
        dff2 <= and_out;
        dff3 <= or_out;
    end

    // Output logic using NOR gate
    assign z = ~(dff1 | dff2 | dff3);

endmodule