module TopModule (
    input logic [2:0] a,
    output logic [15:0] q
);

    always @(*) begin
        case (a)
            3'b000: q = 16'h04D0; // 1232
            3'b001: q = 16'hAEE0; // aee0
            3'b010: q = 16'h27D4; // 27d4
            3'b011: q = 16'h5A0E; // 5a0e
            3'b100: q = 16'h2066; // 2066
            3'b101: q = 16'h64CE; // 64ce
            3'b110: q = 16'hC526; // c526
            3'b111: q = 16'h2F19; // 2f19
            default: q = 16'h0000; // Default case
        endcase
    end

endmodule