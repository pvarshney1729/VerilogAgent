```verilog
module TopModule (
    input logic clk,
    input logic rst, // Added reset input for clarity
    input logic [7:0] in,
    output logic [7:0] anyedge
);

logic [7:0] prev_in; // Internal register to store the previous state of `in`

always @(posedge clk) begin
    if (rst) begin
        anyedge <= 8'b0;
        prev_in <= 8'b0;
    end else begin
        anyedge <= (in ^ prev_in); // XOR operation to detect any edge
        prev_in <= in;
    end
end

endmodule
```