module TopModule (
    output logic out  // 1-bit output, unsigned
);

    // Drive the output to a constant logic low
    assign out = 1'b0;

endmodule