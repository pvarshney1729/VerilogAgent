[BEGIN]
module TopModule (
    input logic [1023:0] in_vector,
    input logic [7:0] select,
    output logic [3:0] out_value
);

    always @(*) begin
        case (select)
            8'd0: out_value = in_vector[3:0];
            8'd1: out_value = in_vector[7:4];
            8'd2: out_value = in_vector[11:8];
            8'd3: out_value = in_vector[15:12];
            8'd4: out_value = in_vector[19:16];
            8'd5: out_value = in_vector[23:20];
            8'd6: out_value = in_vector[27:24];
            8'd7: out_value = in_vector[31:28];
            8'd8: out_value = in_vector[35:32];
            8'd9: out_value = in_vector[39:36];
            8'd10: out_value = in_vector[43:40];
            8'd11: out_value = in_vector[47:44];
            8'd12: out_value = in_vector[51:48];
            8'd13: out_value = in_vector[55:52];
            8'd14: out_value = in_vector[59:56];
            8'd15: out_value = in_vector[63:60];
            8'd16: out_value = in_vector[67:64];
            8'd17: out_value = in_vector[71:68];
            8'd18: out_value = in_vector[75:72];
            8'd19: out_value = in_vector[79:76];
            8'd20: out_value = in_vector[83:80];
            8'd21: out_value = in_vector[87:84];
            8'd22: out_value = in_vector[91:88];
            8'd23: out_value = in_vector[95:92];
            8'd24: out_value = in_vector[99:96];
            8'd25: out_value = in_vector[103:100];
            8'd26: out_value = in_vector[107:104];
            8'd27: out_value = in_vector[111:108];
            8'd28: out_value = in_vector[115:112];
            8'd29: out_value = in_vector[119:116];
            8'd30: out_value = in_vector[123:120];
            8'd31: out_value = in_vector[127:124];
            8'd32: out_value = in_vector[131:128];
            8'd33: out_value = in_vector[135:132];
            8'd34: out_value = in_vector[139:136];
            8'd35: out_value = in_vector[143:140];
            8'd36: out_value = in_vector[147:144];
            8'd37: out_value = in_vector[151:148];
            8'd38: out_value = in_vector[155:152];
            8'd39: out_value = in_vector[159:156];
            8'd40: out_value = in_vector[163:160];
            8'd41: out_value = in_vector[167:164];
            8'd42: out_value = in_vector[171:168];
            8'd43: out_value = in_vector[175:172];
            8'd44: out_value = in_vector[179:176];
            8'd45: out_value = in_vector[183:180];
            8'd46: out_value = in_vector[187:184];
            8'd47: out_value = in_vector[191:188];
            8'd48: out_value = in_vector[195:192];
            8'd49: out_value = in_vector[199:196];
            8'd50: out_value = in_vector[203:200];
            8'd51: out_value = in_vector[207:204];
            8'd52: out_value = in_vector[211:208];
            8'd53: out_value = in_vector[215:212];
            8'd54: out_value = in_vector[219:216];
            8'd55: out_value = in_vector[223:220];
            8'd56: out_value = in_vector[227:224];
            8'd57: out_value = in_vector[231:228];
            8'd58: out_value = in_vector[235:232];
            8'd59: out_value = in_vector[239:236];
            8'd60: out_value = in_vector[243:240];
            8'd61: out_value = in_vector[247:244];
            8'd62: out_value = in_vector[251:248];
            8'd63: out_value = in_vector[255:252];
            8'd64: out_value = in_vector[259:256];
            8'd65: out_value = in_vector[263:260];
            8'd66: out_value = in_vector[267:264];
            8'd67: out_value = in_vector[271:268];
            8'd68: out_value = in_vector[275:272];
            8'd69: out_value = in_vector[279:276];
            8'd70: out_value = in_vector[283:280];
            8'd71: out_value = in_vector[287:284];
            8'd72: out_value = in_vector[291:288];
            8'd73: out_value = in_vector[295:292];
            8'd74: out_value = in_vector[299:296];
            8'd75: out_value = in_vector[303:300];
            8'd76: out_value = in_vector[307:304];
            8'd77: out_value = in_vector[311:308];
            8'd78: out_value = in_vector[315:312];
            8'd79: out_value = in_vector[319:316];
            8'd80: out_value = in_vector[323:320];
            8'd81: out_value = in_vector[327:324];
            8'd82: out_value = in_vector[331:328];
            8'd83: out_value = in_vector[335:332];
            8'd84: out_value = in_vector[339:336];
            8'd85: out_value = in_vector[343:340];
            8'd86: out_value = in_vector[347:344];
            8'd87: out_value = in_vector[351:348];
            8'd88: out_value = in_vector[355:352];
            8'd89: out_value = in_vector[359:356];
            8'd90: out_value = in_vector[363:360];
            8'd91: out_value = in_vector[367:364];
            8'd92: out_value = in_vector[371:368];
            8'd93: out_value = in_vector[375:372];
            8'd94: out_value = in_vector[379:376];
            8'd95: out_value = in_vector[383:380];
            8'd96: out_value = in_vector[387:384];
            8'd97: out_value = in_vector[391:388];
            8'd98: out_value = in_vector[395:392];
            8'd99: out_value = in_vector[399:396];
            8'd100: out_value = in_vector[403:400];
            8'd101: out_value = in_vector[407:404];
            8'd102: out_value = in_vector[411:408];
            8'd103: out_value = in_vector[415:412];
            8'd104: out_value = in_vector[419:416];
            8'd105: out_value = in_vector[423:420];
            8'd106: out_value = in_vector[427:424];
            8'd107: out_value = in_vector[431:428];
            8'd108: out_value = in_vector[435:432];
            8'd109: out_value = in_vector[439:436];
            8'd110: out_value = in_vector[443:440];
            8'd111: out_value = in_vector[447:444];
            8'd112: out_value = in_vector[451:448];
            8'd113: out_value = in_vector[455:452];
            8'd114: out_value = in_vector[459:456];
            8'd115: out_value = in_vector[463:460];
            8'd116: out_value = in_vector[467:464];
            8'd117: out_value = in_vector[471:468];
            8'd118: out_value = in_vector[475:472];
            8'd119: out_value = in_vector[479:476];
            8'd120: out_value = in_vector[483:480];
            8'd121: out_value = in_vector[487:484];
            8'd122: out_value = in_vector[491:488];
            8'd123: out_value = in_vector[495:492];
            8'd124: out_value

// VERILOG-EVAL: response did not use [BEGIN]/[DONE] correctly