```verilog
module TopModule (
    input logic in,  // Input signal
    output logic out // Output signal
);
    assign out = in; // Direct wire behavior
endmodule
```