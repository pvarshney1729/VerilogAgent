module TopModule(
    input logic in,
    output logic out
);
    // Direct wire behavior
    assign out = in;
endmodule