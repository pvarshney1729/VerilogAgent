module TopModule(
    output logic zero
);

// Assign the constant LOW value to the output
assign zero = 1'b0;

endmodule