module TopModule(
    input logic clk,
    input logic resetn,
    input logic x,
    input logic y,
    output logic f,
    output logic g
);

    typedef enum logic [2:0] {
        STATE_A = 3'b000,
        STATE_B = 3'b001,
        STATE_C = 3'b010,
        STATE_D = 3'b011,
        STATE_E = 3'b100,
        STATE_F = 3'b101,
        STATE_G = 3'b110,
        STATE_H = 3'b111
    } state_t;

    state_t current_state, next_state;
    logic [1:0] y_counter;

    // State transition and output logic
    always_ff @(posedge clk) begin
        if (!resetn) begin
            current_state <= STATE_A;
            f <= 0;
            g <= 0;
            y_counter <= 0;
        end else begin
            current_state <= next_state;
            case (current_state)
                STATE_A: begin
                    f <= 0;
                    g <= 0;
                end
                STATE_B: begin
                    f <= 1;
                end
                STATE_C: begin
                    f <= 0;
                end
                STATE_D: begin
                    f <= 0;
                end
                STATE_E: begin
                    f <= 0;
                end
                STATE_F: begin
                    g <= 1;
                end
                STATE_G: begin
                    g <= 1;
                end
                STATE_H: begin
                    g <= 0;
                end
            endcase
        end
    end

    // Next state logic
    always_comb begin
        next_state = current_state;
        case (current_state)
            STATE_A: begin
                if (resetn) next_state = STATE_B;
            end
            STATE_B: begin
                next_state = STATE_C;
            end
            STATE_C: begin
                if (x) next_state = STATE_D;
            end
            STATE_D: begin
                if (!x) next_state = STATE_E;
            end
            STATE_E: begin
                if (x) next_state = STATE_F;
            end
            STATE_F: begin
                if (y) next_state = STATE_G;
                else if (y_counter < 2) y_counter = y_counter + 1;
                else next_state = STATE_H;
            end
            STATE_G: begin
                next_state = STATE_G;
            end
            STATE_H: begin
                next_state = STATE_H;
            end
        endcase
    end

endmodule