module TopModule(
    input  logic in,
    output logic out
);

    // Implement NOT gate logic
    assign out = ~in;

endmodule