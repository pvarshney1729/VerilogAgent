module TopModule
(
  input  logic c,
  input  logic d,
  output logic [3:0] mux_in
);

  // Combinational logic

  assign mux_in[0] = ~c & ~d;
  assign mux_in[1] = c & ~d;
  assign mux_in[2] = c & d;
  assign mux_in[3] = ~c & d;

endmodule