```verilog
module TopModule(
    output logic zero
);
    // Assign constant LOW to the output
    assign zero = 1'b0;
endmodule
```