```verilog
module TopModule (
    input logic clk,  // Clock signal
    input logic ar,   // Asynchronous active-high reset
    input logic d,    // Data input
    output logic q    // D flip-flop output
);
    // D flip-flop implementation with asynchronous reset
    always_ff @(posedge clk or posedge ar) begin
        if (ar) begin
            q <= 1'b0; // Reset output to '0'
        end else begin
            q <= d;    // Capture data input on rising edge of clk
        end
    end
endmodule
```