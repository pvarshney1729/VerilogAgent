module TopModule (
    input logic [3:0] x,
    output logic f
);
    assign f = (x[2] == 1'b0 && x[3] == 1'b0 && (x[0] == 1'b0 && x[1] == 1'b0)) || // 1
                (x[2] == 1'b0 && x[3] == 1'b0 && (x[0] == 1'b1 && x[1] == 1'b0)) || // 0
                (x[2] == 1'b0 && x[3] == 1'b1 && (x[0] == 1'b0 && x[1] == 1'b0)) || // 0
                (x[2] == 1'b0 && x[3] == 1'b1 && (x[0] == 1'b1 && x[1] == 1'b0)) || // 0
                (x[2] == 1'b1 && x[3] == 1'b0 && (x[0] == 1'b0 && x[1] == 1'b0)) || // 1
                (x[2] == 1'b1 && x[3] == 1'b0 && (x[0] == 1'b1 && x[1] == 1'b0)) || // 1
                (x[2] == 1'b1 && x[3] == 1'b1 && (x[0] == 1'b0 && x[1] == 1'b0)) || // 1
                (x[2] == 1'b1 && x[3] == 1'b1 && (x[0] == 1'b1 && x[1] == 1'b0));   // 0
endmodule