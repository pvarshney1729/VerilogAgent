```verilog
module TopModule (
    input logic clk,
    input logic reset,
    input logic in,
    output logic out
);

    typedef enum logic [1:0] {
        A = 2'b00,
        B = 2'b01,
        C = 2'b10,
        D = 2'b11
    } state_t;

    state_t current_state, next_state;

    // State transition logic
    always @(*) begin
        case (current_state)
            A: begin
                if (in) next_state = B;
                else next_state = A;
            end
            B: begin
                if (in) next_state = B;
                else next_state = C;
            end
            C: begin
                if (in) next_state = D;
                else next_state = A;
            end
            D: begin
                if (in) next_state = B;
                else next_state = C;
            end
            default: next_state = A;
        endcase
    end

    // State register and output logic
    always @(posedge clk) begin
        if (reset) begin
            current_state <= A;
            out <= 0;
        end else begin
            current_state <= next_state;
            case (current_state)
                A, B, C: out <= 0;
                D: out <= 1;
                default: out <= 0;
            endcase
        end
    end

endmodule
```