module TopModule (
    input logic clk,        // Clock signal
    input logic reset,      // Synchronous reset signal
    input logic w,          // Control input, 1 bit, unsigned
    output logic Y1,        // Output corresponding to state input y[1]
    output logic Y3         // Output corresponding to state input y[3]
);

    // State encoding
    typedef enum logic [5:0] {
        A = 6'b000001,
        B = 6'b000010,
        C = 6'b000100,
        D = 6'b001000,
        E = 6'b010000,
        F = 6'b100000
    } state_t;

    state_t current_state, next_state;

    // State transition logic
    always @(*) begin
        case (current_state)
            A: next_state = (w) ? B : A;
            B: next_state = (w) ? C : D;
            C: next_state = (w) ? E : D;
            D: next_state = (w) ? F : A;
            E: next_state = (w) ? E : D;
            F: next_state = (w) ? C : D;
            default: next_state = A; // Default to state A for invalid states
        endcase
    end

    // State register with synchronous reset
    always @(posedge clk) begin
        if (reset)
            current_state <= A;
        else
            current_state <= next_state;
    end

    // Output logic
    assign Y1 = current_state[1];
    assign Y3 = current_state[3];

endmodule