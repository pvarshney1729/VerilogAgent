module TopModule(
    input logic in,
    output logic out
);

    // Combinational logic: Direct assignment from input to output
    assign out = in;

endmodule