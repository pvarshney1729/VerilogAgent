```verilog
module TopModule (
    output logic out_one
);

  // Drive the output high continuously
  assign out_one = 1'b1;

endmodule
```