module TopModule(
    output logic zero
);

    // Assign the zero output to logic LOW (0).
    assign zero = 1'b0;

endmodule