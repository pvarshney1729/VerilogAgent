module TopModule(
    output logic out
);

    // Assign a constant logic low (0) to the output 'out'
    assign out = 1'b0;

endmodule