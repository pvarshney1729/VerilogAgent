module TopModule(
    output logic zero
);
    assign zero = 1'b0; // The output is continuously driven to logic LOW (0).
endmodule