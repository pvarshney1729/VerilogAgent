module TopModule(
    output wire out
);
    // Drive the output to logic low
    assign out = 1'b0;
endmodule