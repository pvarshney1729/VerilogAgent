module TopModule (
    input logic clk,
    input logic rst_n,
    input logic [7:0] in,
    output logic [7:0] pedge
);

    logic [7:0] prev_in;

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            prev_in <= 8'b0;
            pedge <= 8'b0;
        end else begin
            pedge <= ~prev_in & in;
            prev_in <= in;
        end
    end

endmodule